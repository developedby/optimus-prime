library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ROM
-- Memoria de programa com 2^15 words de 14 bits

entity rom is
  port (
   clk: in std_logic;
   endereco: in unsigned (14 downto 0);
   dado: out unsigned (13 downto 0)
   );
 end entity;

architecture arq_rom of rom is
  type mem_prog is array (0 to 32767) of unsigned (13 downto 0);
  constant dados_rom : mem_prog := (
        0 => "11000011111111",
        1 => "00000011111001",
        2 => "00111011111001",
        3 => "00011111111001",
        4 => "00000110000011",
        5 => "11000001100100",
        6 => "00000010000100",
        7 => "00000100000000",
        8 => "00100000000011",
        9 => "11111000000001",
        10 => "00000010000011",
        11 => "00000011111000",
        12 => "00000000011000",
        13 => "00001000000100",
        14 => "01110000000000",
        15 => "11001111111001",
        16 => "11000000000001",
        17 => "00000010000011",
        18 => "00100000000011",
        19 => "11111000000001",
        20 => "00000010000011",
        21 => "00000011111000",
        22 => "00000000010000",
        23 => "00100000000010",
        24 => "01100000000000",
        25 => "11001000010001",
        26 => "00000010000101",
        27 => "00000000011001",
        28 => "11000000000001",
        29 => "00001011111001",
        30 => "00100000000101",
        31 => "00000111111000",
        32 => "00001000000100",
        33 => "01110000000001",
        34 => "11001000001000",
        35 => "00011111111000",
        36 => "00000010000110",
        37 => "00000100000000",
        38 => "00000000011000",
        39 => "00100000000110",
        40 => "00011100000101",
        41 => "11001111110111",
        42 => "00100000000011",
        43 => "00001000000100",
        44 => "01110000000000",
        45 => "11001111011111",
    others => (others => '0')
  );
begin
  process(clk)
  begin
    if rising_edge(clk) then
	  dado <= dados_rom(to_integer(endereco));
	end if;
  end process;
end architecture;
